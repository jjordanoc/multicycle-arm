`timescale 1ns/1ps
module controller_tb;

endmodule